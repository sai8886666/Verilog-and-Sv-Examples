// ------------ package --------------

`include "interface.sv"
`include "design1.sv"
`include "transaction.sv"
`include "generator.sv"
`include "coverage.sv"
`include "driver.sv"
`include "input_monitor.sv"
`include "output_monitor.sv"
`include "scorecard.sv"
`include "environment.sv"
`include "test.sv"
`include "top.sv"

