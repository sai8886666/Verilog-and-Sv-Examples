
`include "package.sv"
